module clr_28bit(
    input  wire [27:0] x,
    input  wire [3:0]  y,
    output wire [27:0] r
);

wire d0, d1, t0, t1, t2, t3, t4[27:0], t5[27:0], t6[27:0];

and (t0,y[3],y[0]);
    assign t1 = & {y[2], y[1], t0};
    or (t2,y[1],t0);
        nor (t3,y[2],t2);
            nor (d0,t3,t1);
                not (d1,d0);

assign {t4[27],t4[26],t4[25],t4[24],t4[23],t4[22],t4[21],t4[20],t4[19],t4[18],t4[17],t4[16],t4[15],t4[14],t4[13],t4[12],t4[11],t4[10],t4[9],t4[8],t4[7],t4[6],t4[5],t4[4],t4[3],t4[2],t4[1],t4[0]} =
    {x[26],x[25],x[24],x[23],x[22],x[21],x[20],x[19],x[18],x[17],x[16],x[15],x[14],x[13],x[12],x[11],x[10],x[9],x[8],x[7],x[6],x[5],x[4],x[3],x[2],x[1],x[0],x[27} & {28{d1}};
assign {t5[27],t5[26],t5[25],t5[24],t5[23],t5[22],t5[21],t5[20],t5[19],t5[18],t5[17],t5[16],t5[15],t5[14],t5[13],t5[12],t5[11],t5[10],t5[9],t5[8],t5[7],t5[6],t5[5],t5[4],t5[3],t5[2],t5[1],t5[0]} =
    {x[25],x[24],x[23],x[22],x[21],x[20],x[19],x[18],x[17],x[16],x[15],x[14],x[13],x[12],x[11],x[10],x[9],x[8],x[7],x[6],x[5],x[4],x[3],x[2],x[1],x[0],x[27,x[26]} & {28{d0}};
assign {r[27],r[26],r[25],r[24],r[23],r[22],r[21],r[20],r[19],r[18],r[17],r[16],r[15],r[14],r[13],r[12],r[11],r[10],r[9],r[8],r[7],r[6],r[5],r[4],r[3],r[2],r[1],r[0]} =
    {t4[27],t4[26],t4[25],t4[24],t4[23],t4[22],t4[21],t4[20],t4[19],t4[18],t4[17],t4[16],t4[15],t4[14],t4[13],t4[12],t4[11],t4[10],t4[9],t4[8],t4[7],t4[6],t4[5],t4[4],t4[3],t4[2],t4[1],t4[0]} |
    {t5[27],t5[26],t5[25],t5[24],t5[23],t5[22],t5[21],t5[20],t5[19],t5[18],t5[17],t5[16],t5[15],t5[14],t5[13],t5[12],t5[11],t5[10],t5[9],t5[8],t5[7],t5[6],t5[5],t5[4],t5[3],t5[2],t5[1],t5[0]};

endmodule
