module sbox(
    input  wire [3:0] x,
    output wire [3:0] r
);

wire t0,t1,t2,t3,t4,t5,t6,t7,t8,t9,t10,t11,t12,t13,t14,t15,t16,t17,t18,t19,t20,t21,t22,t23,t24,t25;

not (t0, 3)
not (t1, 2)
and (t2, 2, 0)
nand (t3, 3, 0)
or (t4, 0, 1)
and (t5, 2, 1)
or (t6, 2, 0)
xor (t7, 3, 0)
nor (t8, 2, 1)
xnor (t9, 1, 0)
xor (t10, 3, 2)
    nor (t11, t1, 1)
    and (t12, t6, 3)
    and (t13, t1, 3)
    or (t14, t2, t8)
    nand (t15, t10, t3)
    nand (t16, t2, t0)
    or (t17, t9, t5)
        and (t18, t14, 3)
        nor (t19, t15, 1)
        nor (t20, t12, t2)
        nand (t21, t16, t6)
        and (t22, t13, t4)
        and (t23, t17, t0)
        xor (r[0], t11, t7)
            and (t24, t20, 1)
            and (t25, t21, 1)
            or (r[2], r23, r22)
                or (r[1], t24, t18)
                or (r[2], t25, t19)

endmodule   // 25 gates, 5-gate critical path

/*
Second method, using Karnaugh maps

3210 | r
0000 | 1 1 0 0
0001 | 0 1 0 1
0011 | 1 0 1 1
0010 | 0 1 1 0

0100 | 1 0 0 1
0101 | 0 0 0 0
0111 | 1 1 0 1
0110 | 1 0 1 0

1100 | 0 1 0 0
1101 | 0 1 1 1
1111 | 0 0 1 0
1110 | 0 0 0 1

1000 | 0 0 1 1
1001 | 1 1 1 0
1011 | 1 0 0 0
1010 | 1 1 1 1

r0    32
      00 01 11 10
10 00 0  1  0  1*
   01 1* 0  1* 0
   11 1* 1* 0  0
   10 0  0  1* 1*
0100 | 1101 | 10?0 | 1?10 | 0?11 | 00?1

r1    32
      00 01 11 10
10 00 0  0  0  1*
   01 0  0  1* 1*
   11 1* 0  1* 0
   10 1* 1* 0  1*
0?10 | 001? | 11?1 | 100? | 10?0
0?10 | 001? | 11?1 | 100? | ?010
0?10 | 001? | 11?1 | 1?01 | 10?0

r2    32
      00 01 11 10
10 00 1* 0  1* 0
   01 1* 0  1* 1*
   11 0  1* 0  0
   10 1* 0  0  1*
0111 | ?010 | 110? | 000? | 1?01
0111 | ?010 | 110? | 000? | ?001
0111 | ?010 | 110? | ?001 | 00?0

r3    32
      00 01 11 10
10 00 1* 1* 0  0
   01 0  0  0  1*
   11 1  1  0  1*
   10 0  1  0  1*
10?1 | 101? | 0?00 | 0?11 | 011?
10?1 | 101? | 0?00 | 0?11 | 01?0
10?1 | 101? | 0?00 | 011? | ?011


r0
!3&2&!1&!0 | 3&2&!1&0 | 3&!2&!0 | 3&1&!0 | !3&1&0 | !3&!2&0

r1
!3&1&!0 | !3&!2&1 | 3&2&0 | 3&!2&!1 | 3&!2&!0
!3&1&!0 | !3&!2&1 | 3&2&0 | 3&!2&!1 | !2&1&!0
!3&1&!0 | !3&!2&1 | 3&2&0 | 3&!1&0 | 3&!2&!0

r2
!3&2&1&0 | !2&1&!0 | 3&2&!1 | !3&!2&!1 | 3&!1&0
!3&2&1&0 | !2&1&!0 | 3&2&!1 | !3&!2&!1 | !2&!1&0
!3&2&1&0 | !2&1&!0 | 3&2&!1 | !2&!1&0 | !3&!2&!0

r3
3&!2&0 | 3&!2&1 | !3&!1&!0 | !3&1&0 | !3&2&1
3&!2&0 | 3&!2&1 | !3&!1&!0 | !3&1&0 | !3&2&!0
3&!2&0 | 3&!2&1 | !3&!1&!0 | !3&2&1 | !2&1&0


r0
3^0^(2&!1))
3^0^!(!2 | 1))

r1
1&!(2&0 | 3)        | 3& (2&0 |  !(2 | 0&1))
3& (2&0 | !(2 | 1)) | 1&!(2&0 | 3&(2 | 0))

r2
!1&(!(3^2) | 3&0) | 1&(!3&2&0 | !(2 | 0))
!2&((1^0) | !(3 | 1)) | 2&(!3&1&0 | 3&!1)
!2&((1^0) | !(3 | 0)) | 2&(!3&1&0 | 3&!1)

r3
!3&(!(1^0) | 2&1) | 3&!2&(0 | 1)


t0=!3, t1=!2, t2=2&0, t3=3!&0, t4=0|1, t5=2&1, t6=2|0, t7=3^0, t8=2!|1, t9=1!^0, t10=3^2
t11=t1!|1, t12=t6&3, t13=t1&3, t14=t2|t8, t15=t10!&t3, t16=t2!&t0, t17=t9|t5
t18=t14&3, t19=t15!|1, t20=t12!|t2, t21=t16!&t6, t22=t13&t4, t23=t17&t0
t24=t20&1, t25=t21&1

r0
t11^t7

r1
t24 | t18

r2
t25 | t19

r3
t23 | t22
*/

/*
First method, attempting manual optimisation:
3210 | r
0000 | 1 1 0 0
0001 | 0 1 0 1
0010 | 0 1 1 0
0011 | 1 0 1 1
0100 | 1 0 0 1
0101 | 0 0 0 0
0110 | 1 0 1 0
0111 | 1 1 0 1
1000 | 0 0 1 1
1001 | 1 1 1 0
1010 | 1 1 1 1
1011 | 1 0 0 0
1100 | 0 1 0 0
1101 | 0 1 1 1
1110 | 0 0 0 1
1111 | 0 0 1 0

r0 = 0001 | 0011 | 0100 | 0111 | 1000 | 1010 | 1101 | 1110
r1 = 0010 | 0011 | 0110 | 1000 | 1001 | 1010 | 1101 | 1111
r2 = 0000 | 0001 | 0010 | 0111 | 1001 | 1010 | 1100 | 1101
r3 = 0000 | 0011 | 0100 | 0110 | 0111 | 1001 | 1010 | 1011

r0 = !3&!2&!1&0 | !3&!2&1&0 | !3&2&!1&!0 | !3&2&1&0 | 3&!2&!1&!0 | 3&!2&1&!0 | 3&2&!1&0 | 3&2&1&!0
r1 = !3&!2&1&!0 | !3&!2&1&0 | !3&2&1&!0 | 3&!2&!1&!0 | 3&!2&!1&0 | 3&!2&1&!0 | 3&2&!1&0 | 3&2&1&0
r2 = !3&!2&!1&!0 | !3&!2&!1&0 | !3&!2&1&!0 | !3&2&1&0 | 3&!2&!1&0 | 3&!2&1&!0 | 3&2&!1&!0 | 3&2&!1&0
r3 = !3&!2&!1&!0 | !3&!2&1&0 | !3&2&!1&!0 | !3&2&1&!0 | !3&2&1&0 | 3&!2&!1&0 | 3&!2&1&!0 | 3&!2&1&0

r0 = !3&(!2&0 | 2&!(0^1)) | 3&(!2&!0 | 2&(0^1))
r1 = !3&1&(!2 | 2&!0) | 3&(!2&(!1 | 1&!0) | 2&0)
r2 = !3&(!2&!1 | 1&!(0^2)) | 3&(!2&(0^1) | 2&!1)
r3 = !3&(!2&!(0^1) | 2&(!0 | 1)) | 3&!2&(0 | 1)

r0 = !3&(!2&0 | 2&!(0^1)) | 3&(!(2|0) | 2&(0^1))
r1 = !3&1&!(2&0) | 3&(!(2|1) | !(0^2))
r2 = !3&(!(2|1) | 1&!(0^2)) | 3&(1^(2|0))
r3 = !3&(!(2|(0^1)) | 2&(!0 | 1)) | 3&!2&(0 | 1)

t0=2!|0, t1=1|0, t2=2|1, t3=2&0, t4=!3, t5=0^2, t6=!0, t7=0^1
t9=!t7, t10=!1, t11=2!|t6, t12=2&t9, t13=2&t7, t14=1!^t0, t15=2!|t7, t16=t6|1, t17=t4!|2, t18=t3!|3
t22=t18&1, t23=2&t16, t24=3&t14
t25=t11|t12, t26=t0|t13, t27=t2!&t5, t28=t10|t5, t29=t15|t23, t30=t17&t1
t32=3&t26, t33=3&t27
t34=t4&t25, t35=t22|t33, t36=t2!&t28, t37=t4&t29
t39=t34|t32, t40=t4&t36, t41=t37|t30
t42=t40|t24

r0 = t39
r1 = t35
r2 = t42
r3 = t41

t0=2!|0, t1=1|0, t2=2|1, t3=2&0, t4=!3, t5=0^2, t6=!0, t7=0^1
t8=!t7, t9=!1, t10=2!|t6, t11=2&t8, t12=2&t7, t13=1!^t0, t14=2!|t7, t15=t6|1, t16=t4!|2, t17=t3!|3
t18=t17&1, t19=2&t15, t20=3&t13
t21=t10|t11, t22=t0|t12, t23=t2!&t5, t24=t9|t5, t25=t14|t19, t26=t16&t1
t27=3&t22, t28=3&t23
t29=t4&t21, t30=t18|t28, t31=t2!&t24, t32=t4&t25
t33=t29|t27, t34=t4&t31, t35=t32|t26
t36=t34|t20

r0 = t33
r1 = t30
r2 = t36
r3 = t35


module sbox(
    input  wire [3:0] x,
    output wire [3:0] r
);

wire t0,t1,t2,t3,t4,t5,t6,t7,t8,t9,t10,t11,t12,t13,t14,t15,t16,t17,t18,t19,t20,t21,t22,t23,t24,t25,t26,t27,t28,t29,t30,t31,t32,t33,t34;

nor  (t0, x[2], x[0]);
or   (t1, x[1], x[0]);
or   (t2, x[2], x[1]);
and  (t3, x[2], x[0]);
not  (t4, x[3]);
xor  (t5, x[0], x[2]);
not  (t6, x[0]);
xor  (t7, x[0], x[1]);
not  (t8, x[1]);
xnor (t9, x[0], x[1]);
    nor  (t10, x[2], t6);
    and  (t11, x[2], t9);
    and  (t12, x[2], t7);
    xnor (t13, x[1], t0);
    nor  (t14, x[2], t7);
    or   (t15, x[1], t6);
    nor  (t16, x[2], t4);
    nor  (t17, x[3], t3);
    nand (t23, t2, t5);
    or   (t24, t8, t5);
        and  (t18, x[1], t17);
        and  (t19, x[2], t15);
        and  (t20, x[3], t13);
        or   (t21, t10, t11);
        or   (t22, t0, t12);
        and  (t26, t16, t1);
        and  (t28, x[3], t23);
        nand (t31, t2, t24);
            or   (t25, t14, t19);
            and  (t27, x[3], t22);
            and  (t29, t4, t21);
            or   (r[1], t18, t28);
            and  (t34, t4, t31);
                and  (t32, t4, t25);
                or   (r[0], t29, t27);
                or   (r[2], t34, t20);
                    or   (r[3], t32, t26);

endmodule   // 34 gates, 6-gate critical path
*/